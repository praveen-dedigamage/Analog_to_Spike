** sch_path: /foss/designs/Analog_to_Spike/Schematic/AFE.sch
.subckt AFE

XMsf GND Vin Vsf Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XMb1 Vsf Vb1 Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XC1 Vsf P1 sky130_fd_pr__cap_mim_m3_1 W=16 L=16 m=1
XC2 P1 Vdiff sky130_fd_pr__cap_mim_m3_1 W=4 L=4 m=1
XMr Vdiff Vreset P1 Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XMdp Vdiff P1 Vdd Vdd sky130_fd_pr__pfet_01v8 L=3.2 W=1.5 nf=1 m=1
XMdn Vdiff Vdn GND GND sky130_fd_pr__nfet_01v8 L=3.2 W=1.5 nf=1 m=1
XMONp Vout Vdiff Vdd Vdd sky130_fd_pr__pfet_01v8 L=3.2 W=1.5 nf=1 m=1
XMONn Vout Vonn GND GND sky130_fd_pr__nfet_01v8 L=3.2 W=1.5 nf=1 m=2
Vdd Vdd GND 1.8
vb1 Vb1 GND 0.9
vdn Vdn GND 0.45
voffn Vonn GND 0.5
**** begin user architecture code

** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt




.option savecurrents
.temp 27

* Case #1 -> 100 Hz
Vin vin 0 SIN(0 0.3 100 0 0)
Vreset vreset 0 PULSE(1.8 0 0 1u 1u 900u 1000u)

* Case #2 -> 10 Hz
*Vin vin 0 SIN(0 0.3 10 0 0)
*Vreset vreset 0 PULSE(1.8 0 0 100u 100u 9m 10m)

* Case #3 -> 1 Hz
*Vin vin 0 SIN(0 0.3 1 0 0)
*Vreset vreset 0 PULSE(1.8 0 0 1m 1m 90m 100m)

.control
save all

*Case #1 -> Run 40 ms
tran 1u 0.04

* Case #2 -> Run 400 ms
*tran 100u 0.4

* Case #3 -> Run 4 s
*tran 1m 4


plot vin vout

.endc

**** end user architecture code
.ends
.GLOBAL GND
